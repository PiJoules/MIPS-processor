------------------------------------------------------
-- Adder component
-- Take a wild guess what this does.
------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity adder is
	
end entity;